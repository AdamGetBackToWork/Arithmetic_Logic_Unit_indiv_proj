`ifndef ALU_DEFINES
`define ALU_DEFINES

`define OPER_BITS	2
`define ALU_SUB		`OPER_BITS'b00
`define ALU_LESS	`OPER_BITS'b01
`define ALU_INDB	`OPER_BITS'b10
`define ALU_CHANGE	`OPER_BITS'b11

`endif
