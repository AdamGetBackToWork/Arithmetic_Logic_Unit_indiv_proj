module arith_unit_4

end module
